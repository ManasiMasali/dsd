`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:04:54 03/09/2024 
// Design Name: 
// Module Name:    bcdtoxs3 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bcdtoxs3(b,e);
    input [3:0]b;
    output [3:0]e;
	 assign e[3]=
	 assign e[2]=
	 assign e[1]=
	 assign e[0]=

endmodule
